/*

MIT License

Copyright (c) 2021 7Hemanth

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all
copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
SOFTWARE.

*/

module apb_int(PENABLE,PWRITE,PSEL,PADDR,PWDATA,PRDATA,HWDATA,HRDATA);

input PENABLE,PWRITE;
input [2:0]PSEL;
input [31:0]PADDR,PRDATA,HWDATA;
output reg [31:0]PWDATA,HRDATA;


always@(*) 
begin
	if(PWRITE)
	begin
		if(~PENABLE )
			PWDATA=HWDATA;
		else
			PWDATA=32'bx;
	end
	else if(~PWRITE)
	begin
		if(PENABLE)
			HRDATA=PRDATA;
		else
			HRDATA=32'bx;
	end


end
endmodule